module IF(
  input wire clk,
  input wire i_PC,

  output wire o_PC,
  output wire[31:0] o_imem,
  output wire[31:0] o_inc_pc
  );
endmodule
