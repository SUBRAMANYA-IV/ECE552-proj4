module MEM(
  input wire i_MemWrite,
  input wire[31:0] i_result,
  input wire[31:0] i_address,

  );

endmodule
