module EX(

  );
endmodule
